** Profile: "SCHEMATIC1-trans1"  [ C:\Users\arvba41\OneDrive - Link�pings universitet\Courses\Simulation Course\ODE_Extra_task\battery_task\SPICE\battery_2_state-PSpiceFiles\Voltage_input\battery_2_state_voltage-PSpiceFiles\SCHEMATIC1\trans1.sim ] 

** Creating circuit file "trans1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\arvba41\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3600 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
